package genius_pkg;
    typedef enum logic [1:0] {
        COLOR_RED    = 2'b00,
        COLOR_GREEN  = 2'b01,
        COLOR_BLUE   = 2'b10,
        COLOR_YELLOW = 2'b11
    } color_t;
endpackage